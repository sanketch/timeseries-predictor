module mfdfa(
  input Clk,
  input Rst,
);

  reg [31:0] stocks [300:0] = {107.68, 105.19, 105.67, 106.13, 106.72, 105.91, 105.92, 105.8, 105.97, 104.58, 102.52, 102.26, 101.17, 101.12, 101.03, 101.87, 103.01, 101.5, 100.75, 100.53, 96.69, 96.91, 96.76, 96.1, 94.69, 96.88, 96.04, 96.26, 98.12, 96.64, 93.99, 93.7, 94.27, 94.99, 95.01, 94.02, 96.6, 96.35, 94.48, 96.43, 97.34, 94.09, 93.42, 99.99, 99.44, 101.42, 96.3, 96.79, 96.66, 97.13, 99.52, 97.39, 99.96, 98.53, 96.96, 96.45, 100.7, 102.71, 105.35, 105.26, 107.32, 108.74, 106.82, 108.03, 108.61, 107.23, 107.33, 106.03, 108.98, 111.34, 110.49, 112.48, 113.18, 116.17, 115.62, 118.23, 118.28, 119.03, 115.2, 116.28, 117.34, 118.3, 117.81, 118.03, 118.88, 117.75, 119.3, 118.78, 117.29, 113.69, 114.175, 112.34, 115.72, 116.11, 116.77, 120.57, 121.06, 120.92, 122, 122.57, 121.18, 119.5, 120.53, 119.27, 114.55, 115.28, 119.08, 115.5, 113.76, 113.77, 111.73, 111.04, 111.86, 110.21, 111.79, 111.6, 112.12, 109.5, 110.78, 111.31, 110.78, 110.38, 109.58, 110.3, 109.06, 112.44, 114.71, 115, 114.32, 113.4, 115.21, 113.45, 113.92, 116.41, 116.28, 115.31, 114.21, 112.57, 110.15, 112.31, 109.27, 110.37, 112.34, 107.72, 112.76, 113.29, 112.92, 109.69, 103.74, 103.12, 105.76, 112.65, 115.01, 116.5, 117.16, 115.96, 115.15, 115.24, 113.49, 119.72, 115.52, 115.13, 115.4, 114.64, 118.44, 121.3, 122.37, 122.99, 123.38, 122.77, 124.5, 125.16, 125.22, 130.75, 132.07, 129.62, 128.51, 126.82, 125.61, 125.66, 123.28, 120.07, 122.57, 125.69, 126, 126.44, 126.6, 125.425, 124.53, 126.75, 127.5, 128.11, 127.03, 127.61, 126.6, 127.88, 127.3, 127.6, 126.92, 127.17, 128.59, 128.88, 127.42, 127.8, 128.65, 129.36, 130.12, 129.96, 130.535, 130.28, 131.78, 132.045, 129.62, 132.54, 131.39, 130.06, 130.07, 130.19, 128.77, 128.95, 126.01, 125.865, 126.32, 127.62, 125.26, 125.01, 125.8, 128.7, 128.95, 125.15, 128.64, 130.56, 132.65, 130.28, 129.67, 128.62, 126.91, 127.6, 124.75, 126.17, 126.78, 126.3, 126.85, 127.1, 126.56, 125.6, 126.01, 127.35, 125.32, 124.25, 124.43, 126.37, 123.25, 124.24, 123.38, 126.69, 127.21, 125.9, 127.495, 128.47, 127.04, 124.95, 123.59, 124.45, 122.24, 124.51, 127.14, 126.6, 126.41, 128.54, 129.36, 129.09, 128.46, 130.415, 128.79, 132.17, 133, 129.495, 128.45, 128.715, 127.83, 127.08, 126.46, 124.88, 122.02, 119.72, 118.93, 119.94, 119.56, 118.65, 118.63, 117.16, 118.9, 115.31, 109.14, 113.1, 112.98, 112.4, 109.55, 108.72, 105.99};

parameter MEAN_CALC;
parameter PROFILE_CONSTRUCTION;
parameter CHUNKING;
parameter LOG_RESULTS;


endmodule
